`timescale 1ns / 1ps

module VGA_Syncher (
    input  logic       clk,
    input  logic       reset,
    output logic       h_sync,
    output logic       v_sync,
    output logic       DE,
    output logic [9:0] x_pixel,
    output logic [9:0] y_pixel
);

    logic [9:0] h_counter;
    logic [9:0] v_counter;

    pixel_counter U_Pixel_Counter (.*);
    vgaDecoder U_VGA_Decoder (.*);
endmodule

module pixel_counter (
    input  logic       clk,
    input  logic       reset,
    output logic [9:0] h_counter,
    output logic [9:0] v_counter
);
    localparam H_MAX = 800, V_MAX = 525;

    always_ff @(posedge clk, posedge reset) begin
        if (reset) begin
            h_counter <= 0;
        end else begin
            if (h_counter == H_MAX - 1) begin
                h_counter <= 0;
            end else begin
                h_counter <= h_counter + 1;
            end
        end
    end

    always_ff @(posedge clk, posedge reset) begin
        if (reset) begin
            v_counter <= 0;
        end else begin
            if (h_counter == H_MAX - 1) begin
                if (v_counter == V_MAX - 1) begin
                    v_counter <= 0;
                end else begin
                    v_counter <= v_counter + 1;
                end
            end
        end
    end
endmodule

// module vgaDecoder (
//     input  logic [9:0] h_counter,
//     input  logic [9:0] v_counter,
//     output logic       h_sync,
//     output logic       v_sync,
//     output logic       DE,
//     output logic [9:0] x_pixel,
//     output logic [9:0] y_pixel
// );

    // localparam H_Visible_area = 640;
    // localparam H_Front_porch = 16;
    // localparam H_Sync_pulse = 96;
    // localparam H_Back_porch = 48;

    // localparam V_Visible_area = 480;
    // localparam V_Front_porch = 10;
    // localparam V_Sync_pulse = 2;
    // localparam V_Back_porch = 33;


//     //assign h_sync = !((h_counter >= 656) && (h_counter < 752));
//     assign h_sync = !((h_counter >= H_Visible_area + H_Front_porch) && (h_counter < H_Visible_area + H_Front_porch + H_Sync_pulse));
//     assign v_sync = !((v_counter >= V_Visible_area + V_Front_porch) && (v_counter < V_Visible_area + V_Front_porch + V_Sync_pulse));
//     assign DE = (h_counter < H_Visible_area) && (v_counter < V_Visible_area);
//     assign x_pixel = h_counter;
//     assign y_pixel = v_counter;

// endmodule

module vgaDecoder (
    input  logic       clk,
    input  logic       reset,
    input  logic [9:0] h_counter,
    input  logic [9:0] v_counter,

    output logic       h_sync,
    output logic       v_sync,

    output logic       DE,
    output logic [9:0] x_pixel,
    output logic [9:0] y_pixel
);
    localparam H_Visible_area = 640;
    localparam H_Front_porch  = 16;
    localparam H_Sync_pulse   = 96;

    localparam V_Visible_area = 480;
    localparam V_Front_porch  = 10;
    localparam V_Sync_pulse   = 2;

    // 주소요청용 좌표/DE는 "즉시"
    assign x_pixel = h_counter;
    assign y_pixel = v_counter;
    assign DE      = (h_counter < H_Visible_area) && (v_counter < V_Visible_area);

    // Sync는 comb 계산 후 1clk 지연
    logic h_sync_comb, v_sync_comb;
    assign h_sync_comb =
        !((h_counter >= H_Visible_area + H_Front_porch) &&
          (h_counter <  H_Visible_area + H_Front_porch + H_Sync_pulse));

    assign v_sync_comb =
        !((v_counter >= V_Visible_area + V_Front_porch) &&
          (v_counter <  V_Visible_area + V_Front_porch + V_Sync_pulse));

    always_ff @(posedge clk or posedge reset) begin
        if (reset) begin
            h_sync <= 1'b1;
            v_sync <= 1'b1;
        end else begin
            h_sync <= h_sync_comb;
            v_sync <= v_sync_comb;
        end
    end
endmodule